module regfile(
		input logic clk, we3,
		input logic [4:0] ra1, ra2, wa3,
		input logic [63:0] wd3,
		output logic [63:0] rd1, rd2
	);


	
/* 	logic [63:0] [31:0] registros;
	initial begin
		registros = 32{64'0};
	end
	





	// Leer registros
	always_comb begin

	end */


	// Escribir registros


endmodule