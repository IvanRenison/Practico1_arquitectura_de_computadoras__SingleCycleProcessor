module signext(input logic [31:0] a, output logic [63:0] b);



endmodule
